`timescale 1ns/1ps
module bus_devre (
 input logic [7:0] a,
 output logic [3:0] y
);
assign y = (a == 8'b10000000) ? (4'b0001):
(a == 8'b01000000) ? (4'b0011):
(a==8'b00100000) ? (4'b0010) :
(a== 8'b00010000) ? (4'b0110) :
(a == 8'b00001000) ? (4'b0111) :
(a == 8'b00000100) ? (4'b0101) :
(a ==8'b00000010) ? (4'b0100) :
(a == 8'b00000001)?(4'b1100):(4'b0000);
endmodule
