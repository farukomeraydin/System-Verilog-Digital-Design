`timescale 1ns/1ps
module tb_bus_devre ();
//Bağlanacak giriş-çıkışlar
 logic [7:0] a;
 logic [3:0] y;
// test edeceğimiz devreyi bağlayalım
bus_devre dut0(a,y);
 initial begin
a[7]= 1;a[6] = 0;a[5] = 0; a[4] = 0;a[3] = 0;a[2] = 0;a[1] = 0;a[0] = 0;
#10; //0001
a[7]= 0;a[6] = 1;a[5] = 0; a[4] = 0;a[3] = 0;a[2] = 0;a[1] = 0;a[0] = 0;
#10; //0011
a[7]= 0;a[6] = 0;a[5] = 1; a[4] = 0;a[3] = 0;a[2] = 0;a[1] = 0;a[0] = 0;
#10; //0010
a[7]= 0;a[6] = 0;a[5] = 0; a[4] = 1;a[3] = 0;a[2] = 0;a[1] = 0;a[0] = 0;
#10; //0110
a[7]= 0;a[6] = 0;a[5] = 0; a[4] = 0;a[3] = 1;a[2] = 0;a[1] = 0;a[0] = 0;
#10; //0111
a[7]= 0;a[6] = 0;a[5] = 0; a[4] = 0;a[3] = 0;a[2] = 1;a[1] = 0;a[0] = 0;
#10; //0101
a[7]= 0;a[6] = 0;a[5] = 0; a[4] = 0;a[3] = 0;a[2] = 0;a[1] = 1;a[0] = 0;
#10; //0100
a[7]= 0;a[6] = 0;a[5] = 0; a[4] = 0;a[3] = 0;a[2] = 0;a[1] = 0;a[0] = 1;
#10; //1100
 $stop;
 end
endmodule
